`timescale 1ns / 1ps

module _and(
    input a,
    input b,
    output c
    );
	assign c = a & b;

endmodule
